.circuit
V1 1 GND dc 10    # There can be comment here
I1 GND 1 dc 10
.end
