.circuit
V1 n1 GND ac 5
R2 n1 n2 5
R1 n2 GND 0
.end
