.circuit
I5 1 GND dc 4
I2 GND 2 dc 2
R2 GND 1 2
R6 2 GND 6
R12 2 1 12
.end
